module top(a, sel, out);
  input  [2:0] a;
  input        sel;
  output [1:0] out;
  wire [2:0] a;
  wire       sel;
  wire [1:0] out;
  wire [3:0] z;
  wire w1, w2, w3, w4, w5, \w6 , \1'b1 ,w8;
    not g1 (z[0], a[0]);
    xnor g2 (z[1], a[0], a[1]);
    or g3 (w1, a[0], a[1]);
    xnor g4 (z[2], a[2], w1);
    and g5 (w2, a[2], a[1]);
    and g6 (w3, a[2], a[0]);
    nor g7 (z[3], w2, w3);
    nor g8 (w4, sel, z[3]);
    nor g9 (w5, sel, z[2], 1'b0);
    and g10 ( \w6 , sel, z[1], 1'b1);
    and g11 ( \1'b1 , sel, z[0]);
    or g12 (out[1], w4, \w6 );
    or g13 (out[0], w5, \1'b1 );
endmodule
